// // Copyright (c) 2011-2023 Columbia University, System Level Design Group
// // SPDC-License-Identifier: Apache-2.0

// `timescale 1ps / 1ps
// `include "cache_consts.svh" 
// `include "cache_types.svh" 
// `include "llc_fifo_packet.svh"

// // llc_addr_table.sv 
// // Author: Kevin Jiang
// // processes available incoming signals with priority 

// module llc_addr_table(
//     input llc_addr_t 
// );

// endmodule